LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE work.components.all;

ENTITY Execute IS
--	GENERIC(
--	);
--	PORT(
--	);
END Execute;


ARCHITECTURE structure OF Execute IS
--	signal
BEGIN
END structure;

